module andgate();
